library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Pacote para declarar tipos customizados que serão usados no projeto
package tipos_pacote is
    -- Define um tipo "t_integer_array" como um vetor de inteiros
    type t_integer_array is array (natural range <>) of integer;
end package tipos_pacote;
